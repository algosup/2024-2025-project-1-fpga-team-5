module player (
    output reg [9:0] player_x,
    output reg [9:0] player_y
);

initial begin
    player_x = 10;
    player_y = 15;
end

// Additional logic for player module can  go here

endmodule